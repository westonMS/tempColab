
module example(
    input logic [7:0] sw,
    input logic btnc,
    output logic [3:0] led
);




endmodule